// SPDX-License-Identifier: ISC
`default_nettype none

module cosine (
    input wire clk,
    input  wire [7:0] cos_index,
    output wire [7:0] cos_value,
    output wire zero_pwm
);
  reg zero_pwm_r;
  assign zero_pwm = zero_pwm_r;
  always @(posedge clk) zero_pwm_r <= cos_r == 1'b0;

  reg [7:0] cos_r;
  assign cos_value = cos_r;
  always @(posedge clk)
    case (cos_index)
      8'd0 : cos_r <= 8'd255;
      8'd1 : cos_r <= 8'd255;
      8'd2 : cos_r <= 8'd255;
      8'd3 : cos_r <= 8'd254;
      8'd4 : cos_r <= 8'd254;
      8'd5 : cos_r <= 8'd253;
      8'd6 : cos_r <= 8'd252;
      8'd7 : cos_r <= 8'd251;
      8'd8 : cos_r <= 8'd250;
      8'd9 : cos_r <= 8'd249;
      8'd10 : cos_r <= 8'd247;
      8'd11 : cos_r <= 8'd246;
      8'd12 : cos_r <= 8'd244;
      8'd13 : cos_r <= 8'd242;
      8'd14 : cos_r <= 8'd240;
      8'd15 : cos_r <= 8'd238;
      8'd16 : cos_r <= 8'd236;
      8'd17 : cos_r <= 8'd233;
      8'd18 : cos_r <= 8'd231;
      8'd19 : cos_r <= 8'd228;
      8'd20 : cos_r <= 8'd225;
      8'd21 : cos_r <= 8'd222;
      8'd22 : cos_r <= 8'd219;
      8'd23 : cos_r <= 8'd215;
      8'd24 : cos_r <= 8'd212;
      8'd25 : cos_r <= 8'd208;
      8'd26 : cos_r <= 8'd205;
      8'd27 : cos_r <= 8'd201;
      8'd28 : cos_r <= 8'd197;
      8'd29 : cos_r <= 8'd193;
      8'd30 : cos_r <= 8'd189;
      8'd31 : cos_r <= 8'd185;
      8'd32 : cos_r <= 8'd180;
      8'd33 : cos_r <= 8'd176;
      8'd34 : cos_r <= 8'd171;
      8'd35 : cos_r <= 8'd167;
      8'd36 : cos_r <= 8'd162;
      8'd37 : cos_r <= 8'd157;
      8'd38 : cos_r <= 8'd152;
      8'd39 : cos_r <= 8'd147;
      8'd40 : cos_r <= 8'd142;
      8'd41 : cos_r <= 8'd136;
      8'd42 : cos_r <= 8'd131;
      8'd43 : cos_r <= 8'd126;
      8'd44 : cos_r <= 8'd120;
      8'd45 : cos_r <= 8'd115;
      8'd46 : cos_r <= 8'd109;
      8'd47 : cos_r <= 8'd103;
      8'd48 : cos_r <= 8'd98;
      8'd49 : cos_r <= 8'd92;
      8'd50 : cos_r <= 8'd86;
      8'd51 : cos_r <= 8'd80;
      8'd52 : cos_r <= 8'd74;
      8'd53 : cos_r <= 8'd68;
      8'd54 : cos_r <= 8'd62;
      8'd55 : cos_r <= 8'd56;
      8'd56 : cos_r <= 8'd50;
      8'd57 : cos_r <= 8'd44;
      8'd58 : cos_r <= 8'd37;
      8'd59 : cos_r <= 8'd31;
      8'd60 : cos_r <= 8'd25;
      8'd61 : cos_r <= 8'd19;
      8'd62 : cos_r <= 8'd13;
      8'd63 : cos_r <= 8'd6;
      8'd64 : cos_r <= 8'd0;
      8'd65 : cos_r <= 8'd6;
      8'd66 : cos_r <= 8'd13;
      8'd67 : cos_r <= 8'd19;
      8'd68 : cos_r <= 8'd25;
      8'd69 : cos_r <= 8'd31;
      8'd70 : cos_r <= 8'd37;
      8'd71 : cos_r <= 8'd44;
      8'd72 : cos_r <= 8'd50;
      8'd73 : cos_r <= 8'd56;
      8'd74 : cos_r <= 8'd62;
      8'd75 : cos_r <= 8'd68;
      8'd76 : cos_r <= 8'd74;
      8'd77 : cos_r <= 8'd80;
      8'd78 : cos_r <= 8'd86;
      8'd79 : cos_r <= 8'd92;
      8'd80 : cos_r <= 8'd98;
      8'd81 : cos_r <= 8'd103;
      8'd82 : cos_r <= 8'd109;
      8'd83 : cos_r <= 8'd115;
      8'd84 : cos_r <= 8'd120;
      8'd85 : cos_r <= 8'd126;
      8'd86 : cos_r <= 8'd131;
      8'd87 : cos_r <= 8'd136;
      8'd88 : cos_r <= 8'd142;
      8'd89 : cos_r <= 8'd147;
      8'd90 : cos_r <= 8'd152;
      8'd91 : cos_r <= 8'd157;
      8'd92 : cos_r <= 8'd162;
      8'd93 : cos_r <= 8'd167;
      8'd94 : cos_r <= 8'd171;
      8'd95 : cos_r <= 8'd176;
      8'd96 : cos_r <= 8'd180;
      8'd97 : cos_r <= 8'd185;
      8'd98 : cos_r <= 8'd189;
      8'd99 : cos_r <= 8'd193;
      8'd100 : cos_r <= 8'd197;
      8'd101 : cos_r <= 8'd201;
      8'd102 : cos_r <= 8'd205;
      8'd103 : cos_r <= 8'd208;
      8'd104 : cos_r <= 8'd212;
      8'd105 : cos_r <= 8'd215;
      8'd106 : cos_r <= 8'd219;
      8'd107 : cos_r <= 8'd222;
      8'd108 : cos_r <= 8'd225;
      8'd109 : cos_r <= 8'd228;
      8'd110 : cos_r <= 8'd231;
      8'd111 : cos_r <= 8'd233;
      8'd112 : cos_r <= 8'd236;
      8'd113 : cos_r <= 8'd238;
      8'd114 : cos_r <= 8'd240;
      8'd115 : cos_r <= 8'd242;
      8'd116 : cos_r <= 8'd244;
      8'd117 : cos_r <= 8'd246;
      8'd118 : cos_r <= 8'd247;
      8'd119 : cos_r <= 8'd249;
      8'd120 : cos_r <= 8'd250;
      8'd121 : cos_r <= 8'd251;
      8'd122 : cos_r <= 8'd252;
      8'd123 : cos_r <= 8'd253;
      8'd124 : cos_r <= 8'd254;
      8'd125 : cos_r <= 8'd254;
      8'd126 : cos_r <= 8'd255;
      8'd127 : cos_r <= 8'd255;
      8'd128 : cos_r <= 8'd255;
      8'd129 : cos_r <= 8'd255;
      8'd130 : cos_r <= 8'd255;
      8'd131 : cos_r <= 8'd254;
      8'd132 : cos_r <= 8'd254;
      8'd133 : cos_r <= 8'd253;
      8'd134 : cos_r <= 8'd252;
      8'd135 : cos_r <= 8'd251;
      8'd136 : cos_r <= 8'd250;
      8'd137 : cos_r <= 8'd249;
      8'd138 : cos_r <= 8'd247;
      8'd139 : cos_r <= 8'd246;
      8'd140 : cos_r <= 8'd244;
      8'd141 : cos_r <= 8'd242;
      8'd142 : cos_r <= 8'd240;
      8'd143 : cos_r <= 8'd238;
      8'd144 : cos_r <= 8'd236;
      8'd145 : cos_r <= 8'd233;
      8'd146 : cos_r <= 8'd231;
      8'd147 : cos_r <= 8'd228;
      8'd148 : cos_r <= 8'd225;
      8'd149 : cos_r <= 8'd222;
      8'd150 : cos_r <= 8'd219;
      8'd151 : cos_r <= 8'd215;
      8'd152 : cos_r <= 8'd212;
      8'd153 : cos_r <= 8'd208;
      8'd154 : cos_r <= 8'd205;
      8'd155 : cos_r <= 8'd201;
      8'd156 : cos_r <= 8'd197;
      8'd157 : cos_r <= 8'd193;
      8'd158 : cos_r <= 8'd189;
      8'd159 : cos_r <= 8'd185;
      8'd160 : cos_r <= 8'd180;
      8'd161 : cos_r <= 8'd176;
      8'd162 : cos_r <= 8'd171;
      8'd163 : cos_r <= 8'd167;
      8'd164 : cos_r <= 8'd162;
      8'd165 : cos_r <= 8'd157;
      8'd166 : cos_r <= 8'd152;
      8'd167 : cos_r <= 8'd147;
      8'd168 : cos_r <= 8'd142;
      8'd169 : cos_r <= 8'd136;
      8'd170 : cos_r <= 8'd131;
      8'd171 : cos_r <= 8'd126;
      8'd172 : cos_r <= 8'd120;
      8'd173 : cos_r <= 8'd115;
      8'd174 : cos_r <= 8'd109;
      8'd175 : cos_r <= 8'd103;
      8'd176 : cos_r <= 8'd98;
      8'd177 : cos_r <= 8'd92;
      8'd178 : cos_r <= 8'd86;
      8'd179 : cos_r <= 8'd80;
      8'd180 : cos_r <= 8'd74;
      8'd181 : cos_r <= 8'd68;
      8'd182 : cos_r <= 8'd62;
      8'd183 : cos_r <= 8'd56;
      8'd184 : cos_r <= 8'd50;
      8'd185 : cos_r <= 8'd44;
      8'd186 : cos_r <= 8'd37;
      8'd187 : cos_r <= 8'd31;
      8'd188 : cos_r <= 8'd25;
      8'd189 : cos_r <= 8'd19;
      8'd190 : cos_r <= 8'd13;
      8'd191 : cos_r <= 8'd6;
      8'd192 : cos_r <= 8'd0;
      8'd193 : cos_r <= 8'd6;
      8'd194 : cos_r <= 8'd13;
      8'd195 : cos_r <= 8'd19;
      8'd196 : cos_r <= 8'd25;
      8'd197 : cos_r <= 8'd31;
      8'd198 : cos_r <= 8'd37;
      8'd199 : cos_r <= 8'd44;
      8'd200 : cos_r <= 8'd50;
      8'd201 : cos_r <= 8'd56;
      8'd202 : cos_r <= 8'd62;
      8'd203 : cos_r <= 8'd68;
      8'd204 : cos_r <= 8'd74;
      8'd205 : cos_r <= 8'd80;
      8'd206 : cos_r <= 8'd86;
      8'd207 : cos_r <= 8'd92;
      8'd208 : cos_r <= 8'd98;
      8'd209 : cos_r <= 8'd103;
      8'd210 : cos_r <= 8'd109;
      8'd211 : cos_r <= 8'd115;
      8'd212 : cos_r <= 8'd120;
      8'd213 : cos_r <= 8'd126;
      8'd214 : cos_r <= 8'd131;
      8'd215 : cos_r <= 8'd136;
      8'd216 : cos_r <= 8'd142;
      8'd217 : cos_r <= 8'd147;
      8'd218 : cos_r <= 8'd152;
      8'd219 : cos_r <= 8'd157;
      8'd220 : cos_r <= 8'd162;
      8'd221 : cos_r <= 8'd167;
      8'd222 : cos_r <= 8'd171;
      8'd223 : cos_r <= 8'd176;
      8'd224 : cos_r <= 8'd180;
      8'd225 : cos_r <= 8'd185;
      8'd226 : cos_r <= 8'd189;
      8'd227 : cos_r <= 8'd193;
      8'd228 : cos_r <= 8'd197;
      8'd229 : cos_r <= 8'd201;
      8'd230 : cos_r <= 8'd205;
      8'd231 : cos_r <= 8'd208;
      8'd232 : cos_r <= 8'd212;
      8'd233 : cos_r <= 8'd215;
      8'd234 : cos_r <= 8'd219;
      8'd235 : cos_r <= 8'd222;
      8'd236 : cos_r <= 8'd225;
      8'd237 : cos_r <= 8'd228;
      8'd238 : cos_r <= 8'd231;
      8'd239 : cos_r <= 8'd233;
      8'd240 : cos_r <= 8'd236;
      8'd241 : cos_r <= 8'd238;
      8'd242 : cos_r <= 8'd240;
      8'd243 : cos_r <= 8'd242;
      8'd244 : cos_r <= 8'd244;
      8'd245 : cos_r <= 8'd246;
      8'd246 : cos_r <= 8'd247;
      8'd247 : cos_r <= 8'd249;
      8'd248 : cos_r <= 8'd250;
      8'd249 : cos_r <= 8'd251;
      8'd250 : cos_r <= 8'd252;
      8'd251 : cos_r <= 8'd253;
      8'd252 : cos_r <= 8'd254;
      8'd253 : cos_r <= 8'd254;
      8'd254 : cos_r <= 8'd255;
      default: cos_r <= 8'd255;
    endcase
endmodule
